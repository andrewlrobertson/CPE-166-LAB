module test1(a,b,c);

input a, b;
output c;
and g1(c, a, b);

endmodule